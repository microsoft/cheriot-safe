// Copyright (C) Microsoft Corporation. All rights reserved.




module PULLDOWN ( 
    output O
);

pulldown pd1 (O);

endmodule
