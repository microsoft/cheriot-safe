// Copyright (C) Microsoft Corporation. All rights reserved.




module PULLUP ( 
    output O
);

pullup pd1 (O);

endmodule
